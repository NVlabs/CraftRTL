module stimulus_gen (
        input clk,
        output logic in,
        output logic reset,
        output reg[511:0] wavedrom_title,
        output reg wavedrom_enable,
        input tb_match
);
        task reset_test(input async=0);
                bit arfail, srfail, datafail;

                @(posedge clk);
                @(posedge clk) reset <= 0;
                repeat(3) @(posedge clk);

                @(negedge clk) begin datafail = !tb_match ; reset <= 1; end
                @(posedge clk) arfail = !tb_match;
                @(posedge clk) begin
                        srfail = !tb_match;
                        reset <= 0;
                end
                if (srfail)
                        $display("Hint: Your reset doesn't seem to be working.");
                else if (arfail && (async || !datafail))
                        $display("Hint: Your reset should be %0s, but doesn't appear to be.", async ? "asynchronous" : "synchronous");
                // Don't warn about synchronous reset if the half-cycle before is already wrong. It's more likely
                // a functionality error than the reset being implemented asynchronously.

        endtask


// Add two ports to module stimulus_gen:
//    output [511:0] wavedrom_title
//    output reg wavedrom_enable

        task wavedrom_start(input[511:0] title = "");
        endtask

        task wavedrom_stop;
                #1;
        endtask



        initial begin
                reset <= 1;
                in <= 0;
                @(posedge clk);
                @(posedge clk) reset <= 0; in <= 0;
                @(posedge clk) in <= 1;
                wavedrom_start();
                        // reset_test(0);
                        @(posedge clk) in <= 0;
                        @(posedge clk) in <= 0;
                        @(posedge clk) in <= 0;
                        @(posedge clk) in <= 1;
                        @(posedge clk) in <= 1;
                @(negedge clk);
                wavedrom_stop();
                repeat(30) @(posedge clk, negedge clk) begin
                        in <= $random;
                        // reset <= !($random & 7);
                end

                #1 $finish;
        end

endmodule

module tb();


        wire[511:0] wavedrom_title;
        wire wavedrom_enable;
        int wavedrom_hide_after_time;

        reg clk=0;
        initial forever
                #5 clk = ~clk;

        logic in;
        logic reset;
        logic out;

        initial begin 
                $dumpfile("wave.vcd");
                $dumpvars(1, stim1.clk, clk, reset, in,out );
        end


        wire tb_match;          // Verification
        wire tb_mismatch = ~tb_match;

        stimulus_gen stim1 (
                .clk,
                .* ,
                .in,
                .reset );

        top_module top_module1 (
                .clk,
                .in,
                .reset,
                .out(out) );


        bit strobe = 0;
        task wait_for_end_of_timestep;
                repeat(5) begin
                        strobe <= !strobe;  // Try to delay until the very end of the time step.
                        @(strobe);
                end
        endtask

endmodule